// Digital Design Example
module digital_example (input a, b, output y);
  assign y = a & b;
endmodule
